.param VDD_nom = 5
.param VSS_nom = 0

* Manually step VDD and VSS around nominal (simulate Gaussian samples)
.step param VDD list 4.9 4.91 4.92 4.93 4.94 4.95 4.96 4.97 4.98 4.99 5 5.01 5.02 5.03 5.04 5.05 5.06 5.07 5.08 5.09 5.1
.step param VSS list -0.1 -0.09 -0.08 -0.07 -0.06 -0.05 -0.04 -0.03 -0.02 -0.01 0 0.01 0.02 0.03 0.04 0.05 0.06 0.07 0.08 0.09 0.1

* Voltage sources for Vdd and Vss
Vdd Vdd 0 {VDD}
Vss Vss 0 {VSS}

Vin1 A Vss PULSE(0 {VDD} 0n 10p 10p 10n 20n)
Vin2 B Vss {VDD}

* Load Capacitance
CL Out Vss 1p

* --- NAND Gate (Inverted AND) ---

* PMOS Pull-Up Network (parallel)
M1 NandOut A Vdd Vdd PMOSMOD L=0.18u W=1u
M2 NandOut B Vdd Vdd PMOSMOD L=0.18u W=1u

* NMOS Pull-Down Network (series)
M3 NandOut A Net1 Vss NMOSMOD L=0.18u W=1u
M4 Net1 B Vss Vss NMOSMOD L=0.18u W=1u

* --- Inverter to get final AND Output ---

* PMOS
M5 Out NandOut Vdd Vdd PMOSMOD L=0.18u W=1u

* NMOS
M6 Out NandOut Vss Vss NMOSMOD L=0.18u W=1u

* Default Parameters (fixed now)
.param VTON=0.7
.param VTOP=-0.7
.param KPN=120u
.param KPP=40u

* Models using parameters
.model NMOSMOD NMOS (LEVEL=1 VTO={VTON} KP={KPN})
.model PMOSMOD PMOS (LEVEL=1 VTO={VTOP} KP={KPP})

.tran 0.1n 50n

* --- Delay Measurements Added ---
.meas tran t_rise_in  TRIG V(A) VAL='{VDD}/2' RISE=1 TARG V(A) VAL='{VDD}*0.9' RISE=1
.meas tran t_rise_out TRIG V(Out) VAL='{VDD}/2' RISE=1 TARG V(Out) VAL='{VDD}*0.9' RISE=1
.meas tran delay_param param='t_rise_out - t_rise_in'

.end